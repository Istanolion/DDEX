LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FTOVECT IS
PORT(
	A : IN STD_LOGIC;
	B : IN STD_LOGIC;
	C : IN STD_LOGIC;
	D : IN STD_LOGIC;
	E : IN STD_LOGIC;
	F : IN STD_LOGIC;
	S : OUT STD_LOGIC_VECTOR(0 TO 5)
);
END FTOVECT;

ARCHITECTURE BEHAVORIAL OF FTOVECT IS
	BEGIN
		S(5)<=A;
		S(4)<=B;
		S(3)<=C;
		S(2)<=D;
		S(1)<=E;
		S(0)<=F;
END BEHAVORIAL;