LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FXOR IS
PORT(
	A : IN STD_LOGIC_VECTOR(0 TO 2);
	B : IN STD_LOGIC_VECTOR(0 TO 2);
	S : OUT STD_LOGIC_VECTOR(0 TO 2)
);
END FXOR;

ARCHITECTURE BEHAVORIAL OF FXOR IS
	BEGIN
	S(2)<=A(2) XOR B(2);
	S(1)<=A(1) XOR B(1);
	S(0)<=A(0) XOR B(0);
	END BEHAVORIAL;