LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY NOTF IS
PORT(
	A : IN STD_LOGIC_VECTOR(0 TO 2);
	S : OUT STD_LOGIC_VECTOR(0 TO 2)
);
END NOTF;

ARCHITECTURE BEHAVORIAL OF NOTF IS
	BEGIN
		S(2)<=NOT(A(2));
		S(1)<=NOT(A(1));
		S(0)<=NOT(A(0));
END BEHAVORIAL;