LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MULTPRIN IS
PORT(
	CA2   : IN STD_LOGIC_VECTOR(0 TO 2);
	COMP  : IN STD_LOGIC;
	NOTF  : IN STD_LOGIC_VECTOR(0 TO 2);
	SUMA  : IN STD_LOGIC_VECTOR(0 TO 3);
	RESTA : IN STD_LOGIC_VECTOR(0 TO 3);
	FAND  : IN STD_LOGIC_VECTOR(0 TO 2);
	FXOR  : IN STD_LOGIC_VECTOR(0 TO 2);
	MULT  : IN STD_LOGIC_VECTOR(0 TO 5);
	SELEC : IN STD_LOGIC_VECTOR(0 TO 2);
	S : OUT STD_LOGIC_VECTOR(0 TO 5)
);
END MULTPRIN;

ARCHITECTURE BEHAVORIAL OF MULTPRIN IS
BEGIN
	PROCESS(CA2,COMP,NOTF,SUMA,RESTA,FAND,FXOR,MULT,SELEC)
	BEGIN
		IF (SELEC="000") THEN
			S(5)<=SUMA(3);
			S(4)<=SUMA(2);
			S(3)<=SUMA(1);
			S(2)<=SUMA(0);
			S(1)<='0';
			S(0)<='0';
		ELSIF (SELEC="001") THEN
			S(5)<=RESTA(3);
			S(4)<=RESTA(2);
			S(3)<=RESTA(1);
			S(2)<=RESTA(0);
			S(1)<='0';
			S(0)<='0';
		ELSIF (SELEC="010") THEN
			S(5)<=FAND(2);
			S(4)<=FAND(1);
			S(3)<=FAND(0);
			S(2)<='0';
			S(1)<='0';
			S(0)<='0';
		ELSIF (SELEC="011") THEN
			S(5)<=FXOR(2);
			S(4)<=FXOR(1);
			S(3)<=FXOR(0);
			S(2)<='0';
			S(1)<='0';
			S(0)<='0';
		ELSIF (SELEC="100") THEN
			S(5)<=NOTF(2);
			S(4)<=NOTF(1);
			S(3)<=NOTF(0);
			S(2)<='0';
			S(1)<='0';
			S(0)<='0';
		ELSIF (SELEC="101") THEN
			S(5)<=COMP;
			S(4)<='0';
			S(3)<='0';
			S(2)<='0';
			S(1)<='0';
			S(0)<='0';
		ELSIF (SELEC="110") THEN
			S(5)<=MULT(5);
			S(4)<=MULT(4);
			S(3)<=MULT(3);
			S(2)<=MULT(2);
			S(1)<=MULT(1);
			S(0)<=MULT(0);
		ELSIF (SELEC="111") THEN
			S(5)<=CA2(2);
			S(4)<=CA2(1);
			S(3)<=CA2(0);
			S(2)<='0';
			S(1)<='0';
			S(0)<='0';
		END IF;
	END PROCESS;
END BEHAVORIAL;