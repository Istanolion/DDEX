LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY sUMADOR IS
PORT(
	A : IN STD_LOGIC_VECTOR(0 TO 2);
	B : IN STD_LOGIC_VECTOR(0 TO 2);
	S : OUT STD_LOGIC_VECTOR(0 TO 3)
);
END sUMADOR;

ARCHITECTURE BEHAVORIAL OF SUMADOR IS
	BEGIN
	S(3)<=A(2) XOR B(2);
	S(2)<=(A(2) AND B(2))XOR A(1) XOR B(1);
	S(1)<=(((A(2) AND B(2))AND A(1))  OR  (((A(2) AND B(2))XOR A(1))AND B(1)))XOR A(0) XOR B(0);
	S(0)<=((((A(2) AND B(2))AND A(1))  OR  (((A(2) AND B(2))XOR A(1))AND B(1)))AND A(0))OR(((((A(2) AND B(2))AND A(1))  OR  (((A(2) AND B(2))XOR A(1))AND B(1)))XOR A(0)) AND B(0));   
END BEHAVORIAL;