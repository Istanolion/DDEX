S0<=A0 AND B0;
S1<=(A0 AND B1) XOR(A1 AND B0);
S2<=(A2 AND B0)XOR ((A0 AND B2)XOR(A1 AND B1) XOR ((A1 AND B0) AND (A0 AND B1)));
S3<= (((((A1 AND B0)AND(A0 AND B1))AND((A0 AND B2)XOR(A1 AND B1)))OR((A0 AND B2)AND(A1 AND B1)))XOR((((A1 AND B0)AND(A0 AND B1))XOR((A0 AND B2)XOR(A1 AND B1)))AND(B0 AND A2)))XOR((A1 AND B2)XOR(A2 AND B1));
S4<=()   XOR((((()XOR((((A1 AND B0)AND(A0 AND B1))XOR((A0 AND B2)XOR(A1 AND B1)))AND(A2 AND B0)))AND((A1 AND B2)XOR(A2 AND B1)))OR((A1 AND B2)AND(A2 AND B1)))XOR(A2 AND B2))