LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MUXAB IS 
PORT(
	A : IN STD_LOGIC_VECTOR(0 TO 2);
	B : IN STD_LOGIC_VECTOR(0 TO 2);
	SEL : IN STD_LOGIC;
	OUTPUT : OUT STD_LOGIC_VECTOR(0 TO 2);
	led: out std_logic
);
END MUXAB;

ARCHITECTURE BEHAVIORAL OF MUXAB IS
BEGIN
	PROCESS(A,B,SEL)
	BEGIN
		IF SEL='0' THEN
			OUTPUT<=A;
			led<='1';
		ELSE
			OUTPUT<=B;
			led<='0';
		END IF;
	END PROCESS;
END BEHAVIORAL;