LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY CHANGEBUT IS 
PORT(
	D0 : IN STD_LOGIC;
	OUTPUT : OUT STD_LOGIC
);
END CHANGEBUT;


ARCHITECTURE BEHAVIORAL OF CHANGEBUT IS
SIGNAL SEL: STD_LOGIC:='0';
SIGNAL LASTBUT:STD_LOGIC:='0';
BEGIN
PROCESS(D0)
BEGIN
	IF RISING_EDGE(D0)THEN
	IF(D0='1' AND LASTBUT='0')THEN 
		SEL<=NOT(SEL);
	END IF;
	LASTBUT<=D0;
	OUTPUT<=SEL;
 END IF;
END PROCESS;
END BEHAVIORAL;